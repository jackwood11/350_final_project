module LFSR(NUM_BITS, clk, en, seed, rand_num); 

    input 

endmodule 


  

