module sub_ovf(yes_overflow, A, B, result);
    input [31:0] A, B, result;
    output yes_overflow;

    


endmodule